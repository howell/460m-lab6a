
module microcode_rom(clk, iState, oMicroOp);
    
    input clk;
    input [4:0] iState;
    output [23:0] oMicroOp;

    reg [23:0] rMicrocode [23:0];
    reg [23:0] oMicroOp;

    /* SPR Mux Inputs */
    `define SPR_MUX_INIT        2'd0
    `define SPR_MUX_SPR_SUB_ONE 2'd1
    `define SPR_MUX_SPR_ADD_ONE 2'd2
    
    `define LD_SPR_DIS         1'd0
    `define LD_SPR_EN          1'd1

    /* DAR Mux Select */
    `define DAR_MUX_INIT        2'd0
    `define DAR_MUX_SPR_ADD_ONE 2'd1
    `define DAR_MUX_DAR_SUB_ONE 2'd2
    `define DAR_MUX_DAR_ADD_ONE 2'd3

    `define LD_DAR_DIS          1'd0
    `define LD_DAR_EN           1'd1

    /* DVR Mux Select */
    `define DVR_MUX_INIT    2'd0 
    `define DVR_MUX_DATA_IN 2'd1
    `define DVR_MUX_ALU_OUT 2'd2
    `define DVR_MUX_VAL     2'd3

    `define LD_DVR_DIS      1'd0
    `define LD_DVR_EN       1'd1

    /* Addr Mux Select */
    `define ADDR_MUX_SPR 1'd0
    `define ADDR_MUX_DAR 1'd1

    /* Operand A Mux Select */
    `define OPERAND_A_MUX_DVR     1'd0
    `define OPERAND_A_MUX_DATA_IN 1'd1

    `define LD_OPERAND_A_DIS     1'd0
    `define LD_OPERAND_A_EN      1'd1

    /* Operand B Mux Select */
    `define OPERAND_B_MUX_DVR     1'd0
    `define OPERAND_B_MUX_DATA_IN 1'd1

    `define LD_OPERAND_B_DIS     1'd0
    `define LD_OPERAND_B_EN      1'd1

    /* ALU Select */
    `define ALU_ADD 1'd0
    `define ALU_SUB 1'd1

    /* Data Out Mux */
    `define DATA_OUT_CTRL_MUX_VAL 1'd0
    `define DATA_OUT_CTRL_MUX_ALU 1'd1

    /* Next State Mux Select */
    `define NEXT_STATE_MUX_MICROCODE   1'd0 
    `define NEXT_STATE_MUX_INPUT       1'd1 

    `define CS_DIS          1'd0
    `define CS_EN           1'd1

    `define WE_DIS          1'd0 
    `define WE_EN           1'd1

    `define STATE_PUSH              5'd2
    `define STATE_POP               5'd7
	 `define STATE_ADD               `STATE_ADD_SPR_ADD_ONE_B
	 `define STATE_SUBTRACT          `STATE_SUB_SPR_ADD_ONE_B
	 `define STATE_CLEAR					`STATE_RST
    `define STATE_TOP               `STATE_DAR_SPR_ADD_ONE
	 `define STATE_DEC               `STATE_DEC_DAR
	 `define STATE_INC					`STATE_ADD_DAR
	 
    `define STATE_WAIT              5'd0
    `define STATE_RST               5'd1
    `define STATE_SPR_SPR_SUB_ONE   5'd3 
    `define STATE_DAR_SPR_ADD_ONE   5'd4
    `define STATE_REQUEST_DVR       5'd5
    `define STATE_LOAD_DVR          5'd6
    `define STATE_SUB_SPR_ADD_ONE_B 5'd8
    `define STATE_SUB_REQUEST_B     5'd9
    `define STATE_SUB_LOAD_B        5'd10
    `define STATE_SUB_SPR_ADD_ONE_A 5'd11
    `define STATE_SUB_REQUEST_A     5'd12
    `define STATE_SUB_LOAD_A        5'd13
    `define STATE_SUB_STORE         5'd14
    `define STATE_ADD_SPR_ADD_ONE_B 5'd15
    `define STATE_ADD_REQUEST_B     5'd16
    `define STATE_ADD_LOAD_B        5'd17
    `define STATE_ADD_SPR_ADD_ONE_A 5'd18
    `define STATE_ADD_REQUEST_A     5'd19
    `define STATE_ADD_LOAD_A        5'd20
    `define STATE_ADD_STORE         5'd21
    `define STATE_DEC_DAR           5'd22
    `define STATE_ADD_DAR           5'd23

    initial begin
        rMicrocode[`STATE_WAIT] = {`SPR_MUX_INIT,`LD_SPR_DIS,`DAR_MUX_INIT,
        `LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_INPUT,`CS_DIS,`WE_DIS,`STATE_WAIT};
        rMicrocode[`STATE_RST] = {`SPR_MUX_INIT,`LD_SPR_EN,`DAR_MUX_INIT,
        `LD_DAR_EN,`DVR_MUX_INIT,`LD_DVR_EN,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_WAIT};
        rMicrocode[`STATE_PUSH] = {`SPR_MUX_INIT,`LD_SPR_DIS,`DAR_MUX_INIT,
        `LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_EN,`STATE_SPR_SPR_SUB_ONE};
        rMicrocode[`STATE_SPR_SPR_SUB_ONE] = {`SPR_MUX_SPR_SUB_ONE,
        `LD_SPR_EN,`DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_DAR_SPR_ADD_ONE};
        rMicrocode[`STATE_DAR_SPR_ADD_ONE] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_SPR_ADD_ONE,`LD_DAR_EN,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_REQUEST_DVR};
        rMicrocode[`STATE_REQUEST_DVR] = {`SPR_MUX_INIT,`LD_SPR_DIS,
       `DAR_MUX_SPR_ADD_ONE,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
       `ADDR_MUX_DAR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
       `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
       `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,`STATE_LOAD_DVR};
        rMicrocode[`STATE_LOAD_DVR] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_SPR_ADD_ONE,`LD_DAR_DIS,`DVR_MUX_DATA_IN,`LD_DVR_EN,
        `ADDR_MUX_DAR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,
        `STATE_WAIT};
        rMicrocode[`STATE_POP] = {`SPR_MUX_SPR_ADD_ONE,`LD_SPR_EN,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_DAR_SPR_ADD_ONE};
        rMicrocode[`STATE_SUB_SPR_ADD_ONE_B] = {`SPR_MUX_SPR_ADD_ONE,
        `LD_SPR_EN,`DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_SUB_REQUEST_B};
        rMicrocode[`STATE_SUB_REQUEST_B] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,`STATE_SUB_LOAD_B};
        rMicrocode[`STATE_SUB_LOAD_B] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DATA_IN,
        `LD_OPERAND_B_EN,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_SUB_SPR_ADD_ONE_A};
        rMicrocode[`STATE_SUB_SPR_ADD_ONE_A] = {`SPR_MUX_SPR_ADD_ONE,
        `LD_SPR_EN,`DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_SUB_REQUEST_A};
        rMicrocode[`STATE_SUB_REQUEST_A] ={`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,`STATE_SUB_LOAD_A};
        rMicrocode[`STATE_SUB_LOAD_A] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DATA_IN,`LD_OPERAND_A_EN,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_SUB_STORE};
        rMicrocode[`STATE_SUB_STORE] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_ALU_OUT,`LD_DVR_EN,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_SUB,
        `DATA_OUT_CTRL_MUX_ALU,`NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_EN,
        `STATE_SPR_SPR_SUB_ONE};
        rMicrocode[`STATE_ADD_SPR_ADD_ONE_B] = {`SPR_MUX_SPR_ADD_ONE,
        `LD_SPR_EN,`DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_ADD_REQUEST_B};
        rMicrocode[`STATE_ADD_REQUEST_B] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,`STATE_ADD_LOAD_B};
        rMicrocode[`STATE_ADD_LOAD_B] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DATA_IN,
        `LD_OPERAND_B_EN,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_ADD_SPR_ADD_ONE_A};
        rMicrocode[`STATE_ADD_SPR_ADD_ONE_A] = {`SPR_MUX_SPR_ADD_ONE,
        `LD_SPR_EN,`DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_ADD_REQUEST_A};
        rMicrocode[`STATE_ADD_REQUEST_A] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_DIS,`STATE_ADD_LOAD_A};
        rMicrocode[`STATE_ADD_LOAD_A] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_INIT,`LD_DVR_DIS,`ADDR_MUX_SPR,
        `OPERAND_A_MUX_DATA_IN,`LD_OPERAND_A_EN,`OPERAND_B_MUX_DVR,
        `LD_OPERAND_B_DIS,`ALU_ADD,`DATA_OUT_CTRL_MUX_VAL,
        `NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,`STATE_ADD_STORE};
        rMicrocode[`STATE_ADD_STORE] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_INIT,`LD_DAR_DIS,`DVR_MUX_ALU_OUT,`LD_DVR_EN,
        `ADDR_MUX_SPR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_ALU,`NEXT_STATE_MUX_MICROCODE,`CS_EN,`WE_EN,
        `STATE_SPR_SPR_SUB_ONE};
        rMicrocode[`STATE_DEC_DAR] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_DAR_SUB_ONE,`LD_DAR_EN,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_DAR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_REQUEST_DVR};
        rMicrocode[`STATE_ADD_DAR] = {`SPR_MUX_INIT,`LD_SPR_DIS,
        `DAR_MUX_DAR_ADD_ONE,`LD_DAR_EN,`DVR_MUX_INIT,`LD_DVR_DIS,
        `ADDR_MUX_DAR,`OPERAND_A_MUX_DVR,`LD_OPERAND_A_DIS,
        `OPERAND_B_MUX_DVR,`LD_OPERAND_B_DIS,`ALU_ADD,
        `DATA_OUT_CTRL_MUX_VAL,`NEXT_STATE_MUX_MICROCODE,`CS_DIS,`WE_DIS,
        `STATE_REQUEST_DVR};
    end

    always @(negedge clk) begin
        if(~clk) begin
            oMicroOp <= rMicrocode[iState]; 
        end
        else begin
        end
    end /* always */

endmodule /* microcode_rom */
